/*******************************************************
** NAME: common
** DESC: define some configs
********************************************************/

// Enable ILA
// `define DEBUG


`define PERF_MON